-- megafunction wizard: %RAM: 1-PORT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altsyncram 

-- ============================================================
-- File Name: RAM.vhd
-- Megafunction Name(s):
-- 			altsyncram
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 16.1.2 Build 203 01/18/2017 SJ Standard Edition
-- ************************************************************


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY altera_mf;
USE altera_mf.altera_mf_components.all;

ENTITY RAM IS
	GENERIC(
		DataWidth : INTEGER := 8;
		AddrWidth : INTEGER := 9
	);
	PORT(
		address : IN STD_LOGIC_VECTOR ( ( AddrWidth - 1 ) DOWNTO 0 );
		clock   : IN STD_LOGIC := '1';
		data    : IN STD_LOGIC_VECTOR ( ( DataWidth - 1 ) DOWNTO 0 );
		rden    : IN STD_LOGIC := '1';
		wren    : IN STD_LOGIC;
		q       : OUT STD_LOGIC_VECTOR ( ( DataWidth - 1 ) DOWNTO 0 )
	);
END RAM;


ARCHITECTURE SYN OF ram IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR ( ( DataWidth - 1 ) DOWNTO 0 );

BEGIN
	q    <= sub_wire0( ( DataWidth - 1 ) DOWNTO 0 );

	altsyncram_component : altsyncram
	GENERIC MAP (
		clock_enable_input_a => "BYPASS",
		clock_enable_output_a => "BYPASS",
		intended_device_family => "Cyclone IV GX",
		lpm_hint => "ENABLE_RUNTIME_MOD=NO",
		lpm_type => "altsyncram",
		numwords_a => ( 2 ** AddrWidth ),
		operation_mode => "SINGLE_PORT",
		outdata_aclr_a => "NONE",
		outdata_reg_a => "CLOCK0",
		power_up_uninitialized => "FALSE",
		--read_during_write_mode_port_a => "OLD_DATA",
		widthad_a => AddrWidth,
		width_a => DataWidth,
		width_byteena_a => 1
	)
	PORT MAP (
		address_a => address,
		clock0 => clock,
		data_a => data,
		rden_a => rden,
		wren_a => wren,
		q_a => sub_wire0
	);



END SYN;

