`define hash 32'hf49cd86
`define timestmp 1655817855
`define number_version 2958367
