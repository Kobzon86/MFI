LIBRARY IEEE;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.STD_LOGIC_1164.ALL;

PACKAGE key_codes_pkg IS

	---------- String Select KEYS -----------------
	CONSTANT KEY_LEFT1   : INTEGER := 400;
	CONSTANT KEY_RIGHT1  : INTEGER := 401;
	CONSTANT KEY_LEFT2   : INTEGER := 402;
	CONSTANT KEY_RIGHT2  : INTEGER := 403;
	CONSTANT KEY_LEFT3   : INTEGER := 404;
	CONSTANT KEY_RIGHT3  : INTEGER := 405;	
	CONSTANT KEY_LEFT4   : INTEGER := 406;
	CONSTANT KEY_RIGHT4  : INTEGER := 407;	
	CONSTANT KEY_LEFT5   : INTEGER := 408;
	CONSTANT KEY_RIGHT5  : INTEGER := 409;
	CONSTANT KEY_LEFT6   : INTEGER := 410;
	CONSTANT KEY_RIGHT6  : INTEGER := 411;	
	CONSTANT KEY_LEFT7   : INTEGER := 412;
	CONSTANT KEY_RIGHT7  : INTEGER := 413;
	CONSTANT KEY_LEFT8   : INTEGER := 414;
	CONSTANT KEY_RIGHT8  : INTEGER := 415;
	CONSTANT KEY_LEFT9   : INTEGER := 416;
	CONSTANT KEY_RIGHT9  : INTEGER := 417;
	CONSTANT KEY_LEFT10  : INTEGER := 418;
	CONSTANT KEY_RIGHT10 : INTEGER := 419;
	--------- NEW KEYS MFI2-15 ------------------
	CONSTANT KEY_LEFT11  : INTEGER := 452;
	CONSTANT KEY_RIGHT11 : INTEGER := 453;
	CONSTANT KEY_LEFT12  : INTEGER := 454;
	CONSTANT KEY_RIGHT12 : INTEGER := 455;
	CONSTANT KEY_LEFT13  : INTEGER := 456;
	CONSTANT KEY_RIGHT13 : INTEGER := 457;
	CONSTANT KEY_LEFT14  : INTEGER := 458;
	CONSTANT KEY_RIGHT14 : INTEGER := 459;
	CONSTANT KEY_LEFT15  : INTEGER := 460;
	CONSTANT KEY_RIGHT15 : INTEGER := 461;
	CONSTANT KEY_LEFT16  : INTEGER := 462;
	CONSTANT KEY_RIGHT16 : INTEGER := 463;
	
	
	
	---------- Column Select KEYS -----------------
	CONSTANT KEY_UP1    : INTEGER := 420;
	CONSTANT KEY_DOWN1  : INTEGER := 421;
	CONSTANT KEY_UP2    : INTEGER := 422;
	CONSTANT KEY_DOWN2  : INTEGER := 423;
	CONSTANT KEY_UP3    : INTEGER := 424;
	CONSTANT KEY_DOWN3  : INTEGER := 425;	
	CONSTANT KEY_UP4    : INTEGER := 426;
	CONSTANT KEY_DOWN4  : INTEGER := 427;	
	CONSTANT KEY_UP5    : INTEGER := 428;
	CONSTANT KEY_DOWN5  : INTEGER := 429;
	CONSTANT KEY_UP6    : INTEGER := 430;
	CONSTANT KEY_DOWN6  : INTEGER := 431;	
	CONSTANT KEY_UP7    : INTEGER := 432;
	CONSTANT KEY_DOWN7  : INTEGER := 433;
	CONSTANT KEY_UP8    : INTEGER := 434;
	CONSTANT KEY_DOWN8  : INTEGER := 435;
	CONSTANT KEY_UP9    : INTEGER := 436;
	CONSTANT KEY_DOWN9  : INTEGER := 437;
	CONSTANT KEY_UP10   : INTEGER := 438;
	CONSTANT KEY_DOWN10 : INTEGER := 439;
	--------- NEW KEYS MFI2-15 --------------
	CONSTANT KEY_UP11   : INTEGER := 440;
	CONSTANT KEY_DOWN11 : INTEGER := 441;
	CONSTANT KEY_UP12   : INTEGER := 442;
	CONSTANT KEY_DOWN12 : INTEGER := 443;
	CONSTANT KEY_UP13   : INTEGER := 444;
	CONSTANT KEY_DOWN13 : INTEGER := 445;
	CONSTANT KEY_UP14   : INTEGER := 446;
	CONSTANT KEY_DOWN14 : INTEGER := 447;
	CONSTANT KEY_UP15   : INTEGER := 448;
	CONSTANT KEY_DOWN15 : INTEGER := 449;
	CONSTANT KEY_UP16   : INTEGER := 450;
	CONSTANT KEY_DOWN16 : INTEGER := 451;
	
	


	----------- FUNCTIONAL KEYS -----------------
	CONSTANT KEY_DATA    : INTEGER := 600;
	CONSTANT KEY_NAV     : INTEGER := 601;
	CONSTANT KEY_VNAV    : INTEGER := 602;
	CONSTANT KEY_DTO     : INTEGER := 603;
	CONSTANT KEY_LIST    : INTEGER := 604;
	CONSTANT KEY_PREV    : INTEGER := 605;
	CONSTANT KEY_FUEL    : INTEGER := 606;
	CONSTANT KEY_FPL     : INTEGER := 607;
	CONSTANT KEY_PERF    : INTEGER := 608;
	CONSTANT KEY_TUNE    : INTEGER := 609;
	CONSTANT KEY_MENU    : INTEGER := 610;
	CONSTANT KEY_NEXT    : INTEGER := 611;
	CONSTANT KEY_BACK    : INTEGER := 612;
	CONSTANT KEY_MSG     : INTEGER := 613;
	CONSTANT KEY_CTRL    : INTEGER := 614;
	CONSTANT KEY_ENTER   : INTEGER := 615;
	CONSTANT KEY_SIGN    : INTEGER := 616;
	CONSTANT KEY_ADSB    : INTEGER := 617;
	CONSTANT KEY_ABC     : INTEGER := 619;
	CONSTANT KEY_123     : INTEGER := 620;
	CONSTANT KEY_LEFT    : INTEGER := 621;
	CONSTANT KEY_TAWS    : INTEGER := 622;
	CONSTANT KEY_RIGHT   : INTEGER := 624;
	CONSTANT KEY_SEL     : INTEGER := 625;
	CONSTANT KEY_SLASH   : INTEGER := 626;
	CONSTANT KEY_DOT     : INTEGER := 627;
	CONSTANT KEY_TRFC    : INTEGER := 628;
	CONSTANT KEY_WXR     : INTEGER := 629;
	CONSTANT KEY_MODE    : INTEGER := 630;
	
	
	--------- NUMERIC KEYS ----------------------
	CONSTANT KEY_0       : INTEGER := 548;
	CONSTANT KEY_1       : INTEGER := 549;
	CONSTANT KEY_2       : INTEGER := 550;
	CONSTANT KEY_3       : INTEGER := 551;
	CONSTANT KEY_4       : INTEGER := 552;
	CONSTANT KEY_5       : INTEGER := 553;
	CONSTANT KEY_6       : INTEGER := 554;
	CONSTANT KEY_7       : INTEGER := 555;
	CONSTANT KEY_8       : INTEGER := 556;
	CONSTANT KEY_9       : INTEGER := 557;
	
	----------- ABC KEYS ------------------------
	CONSTANT KEY_A       : INTEGER := 565;
	CONSTANT KEY_B       : INTEGER := 566;
	CONSTANT KEY_C       : INTEGER := 567;
	CONSTANT KEY_D       : INTEGER := 568;
	CONSTANT KEY_E       : INTEGER := 569;
	CONSTANT KEY_F       : INTEGER := 570;
	CONSTANT KEY_G       : INTEGER := 571;
	CONSTANT KEY_H       : INTEGER := 572;
	CONSTANT KEY_I       : INTEGER := 573;
	CONSTANT KEY_J       : INTEGER := 574;
	CONSTANT KEY_K       : INTEGER := 575;
	CONSTANT KEY_L       : INTEGER := 576;
	CONSTANT KEY_M       : INTEGER := 577;
	CONSTANT KEY_N       : INTEGER := 578;
	CONSTANT KEY_O       : INTEGER := 579;
	CONSTANT KEY_P       : INTEGER := 580;
	CONSTANT KEY_Q       : INTEGER := 581;
	CONSTANT KEY_R       : INTEGER := 582;
	CONSTANT KEY_S       : INTEGER := 583;
	CONSTANT KEY_T       : INTEGER := 584;
	CONSTANT KEY_U       : INTEGER := 585;
	CONSTANT KEY_V       : INTEGER := 586;
	CONSTANT KEY_W       : INTEGER := 587;
	CONSTANT KEY_X       : INTEGER := 588;
	CONSTANT KEY_Y       : INTEGER := 589;
	CONSTANT KEY_Z       : INTEGER := 590;
	
	--------- Valcoders Buttons functions assign -------------
	CONSTANT VALLEFT_BTN  : INTEGER := KEY_CTRL; -- VAL1_BTN
	CONSTANT VALRIGHT_BTN : INTEGER := KEY_SEL; -- VAL2_BTN
	
	CONSTANT NO_KEY      : INTEGER := 0;
	
	CONSTANT WORD_0370_CODE_START : INTEGER := KEY_DATA;
	CONSTANT WORD_0370_CODE_STOP  : INTEGER := KEY_ADSB;
	CONSTANT WORD_0371_CODE_START : INTEGER := KEY_ABC;
	CONSTANT WORD_0371_CODE_STOP  : INTEGER := KEY_WXR;
	--CONSTANT WORD_0372_CODE_START : INTEGER := KEY_DATA; --
	--CONSTANT WORD_0372_CODE_STOP  : INTEGER := KEY_ADSB; --
	CONSTANT WORD_0373_CODE_START : INTEGER := KEY_LEFT1; 
	CONSTANT WORD_0373_CODE_STOP  : INTEGER := KEY_RIGHT9; 
	--CONSTANT WORD_0373_CODE_STOP  : INTEGER := KEY_RIGHT10; 
	CONSTANT WORD_0374_CODE_START : INTEGER := KEY_UP1; 
	CONSTANT WORD_0374_CODE_STOP  : INTEGER := KEY_DOWN9;
	--CONSTANT WORD_0374_CODE_STOP  : INTEGER := KEY_DOWN10; 
	
	--CONSTANT WORD_0375_CODE_START : INTEGER := KEY_ABC; --
	--CONSTANT WORD_0375_CODE_STOP  : INTEGER := KEY_WXR; --
	--CONSTANT WORD_0376_CODE_START : INTEGER := KEY_DATA; --
	--CONSTANT WORD_0376_CODE_STOP  : INTEGER := KEY_ADSB; --
	--CONSTANT WORD_0377_CODE_START : INTEGER := KEY_ABC; --
	--CONSTANT WORD_0377_CODE_STOP  : INTEGER := KEY_WXR; --
	
	CONSTANT WORD_0357_CODE_START   : INTEGER := KEY_UP10;
	CONSTANT WORD_0357_CODE_STOP    : INTEGER := KEY_DOWN16;


END key_codes_pkg;
