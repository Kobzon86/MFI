LIBRARY IEEE;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.STD_LOGIC_1164.ALL;


PACKAGE milstd_1553_pkg IS

	CONSTANT FreqMult              : INTEGER := 16;
	CONSTANT RAM_RX_ADDR_WIDTH_PKG : INTEGER := 12; --12;
	CONSTANT RAM_TX_ADDR_WIDTH_PKG : INTEGER := RAM_RX_ADDR_WIDTH_PKG; --12;
	CONSTANT RAM_DATA_WIDTH_PKG    : INTEGER := 32;
	
	---------------- line signals constants -------------------
	CONSTANT SYNC_TYPE_DATA : STD_LOGIC_VECTOR( 1 DOWNTO 0 ) := "01";
	CONSTANT SYNC_TYPE_COMM : STD_LOGIC_VECTOR( 1 DOWNTO 0 ) := "10";
	CONSTANT SYNC_TYPE_PAUSE : STD_LOGIC_VECTOR( 1 DOWNTO 0 ) := "11";
		
	CONSTANT TX_SYNC_DATA   : STD_LOGIC_VECTOR( 11 DOWNTO 0 ) := "000000111111";
	CONSTANT TX_SYNC_COMM   : STD_LOGIC_VECTOR( 11 DOWNTO 0 ) := "111111000000"; --"111110000000"
	
	CONSTANT SYNC_COMSTAT : STD_LOGIC_VECTOR( ( ( FreqMult * 3 ) - 1 ) DOWNTO 0 ) := x"7FFFFF000000"; --x"FFFFFF000000";
	CONSTANT SYNC_COMSTAT2: STD_LOGIC_VECTOR( ( ( FreqMult * 3 ) - 1 ) DOWNTO 0 ) := x"FFFFFF000000"; --x"FFFFFF000000";
	
	CONSTANT SYNC_DATA    : STD_LOGIC_VECTOR( ( ( FreqMult * 3 ) - 1 ) DOWNTO 0 ) := x"0000007FFFFF";
	CONSTANT SYNC_DATA2   : STD_LOGIC_VECTOR( ( ( FreqMult * 3 ) - 1 ) DOWNTO 0 ) := x"8000007FFFFF";
	CONSTANT SYNC_DATA3   : STD_LOGIC_VECTOR( ( ( FreqMult * 3 ) - 1 ) DOWNTO 0 ) := x"8000003FFFFF";
	CONSTANT SYNC_DATA4   : STD_LOGIC_VECTOR( ( ( FreqMult * 3 ) - 1 ) DOWNTO 0 ) := x"0000007FFFFE";	
	
	CONSTANT TX_SYNC_LEN    : UNSIGNED( 7 DOWNTO 0 ) := x"0C"; --x"06";	
	CONSTANT TX_WRD_LEN     : UNSIGNED( 7 DOWNTO 0 ) := x"50";--x"28";	-- 20 bits 
	
	CONSTANT BROAD_ADDR     : STD_LOGIC_VECTOR( 4 DOWNTO 0 ) := "11111";
	CONSTANT DRV_MODE_1     : STD_LOGIC_VECTOR( 4 DOWNTO 0 ) := "11111";
	CONSTANT DRV_MODE_0     : STD_LOGIC_VECTOR( 4 DOWNTO 0 ) := "00000";

	CONSTANT RX_TRANSACT    : STD_LOGIC := '0';
	CONSTANT TX_TRANSACT    : STD_LOGIC := '1';

	---------------- command codes without TxRx bit ---------------------------
	CONSTANT DYN_BUS_CNTL                 : STD_LOGIC_VECTOR( 4 DOWNTO 0 ) := "00000";
	CONSTANT SYNCHRONIZE                  : STD_LOGIC_VECTOR( 4 DOWNTO 0 ) := "00001";
	CONSTANT TX_STAT_WRD                  : STD_LOGIC_VECTOR( 4 DOWNTO 0 ) := "00010";
	CONSTANT INIT_SELFTEST                : STD_LOGIC_VECTOR( 4 DOWNTO 0 ) := "00011";
	CONSTANT TRANS_SHUTDWN                : STD_LOGIC_VECTOR( 4 DOWNTO 0 ) := "00100";
	CONSTANT OVRD_TRANS_SHUTDWN           : STD_LOGIC_VECTOR( 4 DOWNTO 0 ) := "00101"; 
	CONSTANT INHIB_TERMIN_FLAG            : STD_LOGIC_VECTOR( 4 DOWNTO 0 ) := "00110";
	CONSTANT OVRD_INHIB_TERMIN_FLAG       : STD_LOGIC_VECTOR( 4 DOWNTO 0 ) := "00111";
	CONSTANT RST_REMOTE_TERMINAL          : STD_LOGIC_VECTOR( 4 DOWNTO 0 ) := "01000";
	CONSTANT TX_VECTOR_WRD                : STD_LOGIC_VECTOR( 4 DOWNTO 0 ) := "10000";
	CONSTANT SYNCHRONIZE_DWRD             : STD_LOGIC_VECTOR( 4 DOWNTO 0 ) := "10001";
	CONSTANT TX_LAST_COMAND               : STD_LOGIC_VECTOR( 4 DOWNTO 0 ) := "10010";
	CONSTANT TX_BIT_WORD                  : STD_LOGIC_VECTOR( 4 DOWNTO 0 ) := "10011";
	CONSTANT SELECTED_TRANS_SHUTDWN       : STD_LOGIC_VECTOR( 4 DOWNTO 0 ) := "10100";
	CONSTANT OVRD_SELECTED_TRANS_SHUTDWN  : STD_LOGIC_VECTOR( 4 DOWNTO 0 ) := "10101";

	---------------------- RXTX_Buffer settings  --------------------------------
	CONSTANT BUFF_LEN_BYTES   : UNSIGNED( 15 DOWNTO 0 ) := TO_UNSIGNED( 2048, 16 );
	CONSTANT BUFF_LEN_WORDS   : UNSIGNED( 15 DOWNTO 0 ) := TO_UNSIGNED( 512, 16 );
	CONSTANT SECTOR_LEN_WORDS : UNSIGNED( RAM_RX_ADDR_WIDTH_PKG DOWNTO 0 ) := TO_UNSIGNED( 32, RAM_RX_ADDR_WIDTH_PKG + 1 ); -- SECTOR LEN for SubAddress
	
	------------------- REGISTERS addresses ----------------------
	CONSTANT CONFIG_REG_ADDR   : INTEGER := 0;
	CONSTANT INTMASK_REG_ADDR  : INTEGER := 1;
	CONSTANT INTFLAG_REG_ADDR  : INTEGER := 2;
	CONSTANT STATE_REG_ADDR    : INTEGER := 3;
	CONSTANT ADDRMASK_REG_ADDR : INTEGER := 4; 

	----------- CONFIG_REG bits ---------------------
	CONSTANT CPU_BUFF_BUSY : INTEGER := 26; -- Moved from STATE_REG
	CONSTANT SOFT_NODEADDR : INTEGER := 24;
	CONSTANT TST_TXCHANNEL : INTEGER := 23;
	CONSTANT TST_NADDR_H   : INTEGER := 22;
	CONSTANT TST_NADDR_L   : INTEGER := 18;
	CONSTANT TST_SADDR_H   : INTEGER := 17;
	CONSTANT TST_SADDR_L   : INTEGER := 13;
	CONSTANT TST_WRDSNUM_H : INTEGER := 12;
	CONSTANT TST_WRDSNUM_L : INTEGER := 8;
	CONSTANT LINE_OFF      : INTEGER := 7;
	CONSTANT DIAG          : INTEGER := 6;
	CONSTANT RXTX_EN       : INTEGER := 5;
	CONSTANT NODE_ADDR_H   : INTEGER := 4;
	CONSTANT NODE_ADDR_L   : INTEGER := 0;
	
	---------- INTFLAG_REG bits --------------------
	CONSTANT TX_ERROR1     : INTEGER := 3;  -- Moved from STATE_REG
	CONSTANT TX_ERROR2     : INTEGER := 2;  -- Moved from STATE_REG
	CONSTANT TX_COMPL      : INTEGER := 1;
	CONSTANT RX_OK         : INTEGER := 0;
	
	
	---------- STATE_REG bits ----------------------
	CONSTANT HARD_NODEADDR_H : INTEGER := 27; -- MUST BE USED!! but not used yet
	CONSTANT HARD_NODEADDR_L : INTEGER := 23; -- MUST BE USED!! but not used yet
	CONSTANT RXWRD_CNT_H    : INTEGER := 22;
	CONSTANT RXWRD_CNT_L    : INTEGER := 17;
	CONSTANT RX_LASTSUB_H   : INTEGER := 16;
	CONSTANT RX_LASTSUB_L   : INTEGER := 12;
	CONSTANT FPGA_BUFF_BUSY : INTEGER := 8;
	CONSTANT MSG_ERR        : INTEGER := 7;
	CONSTANT INSTR          : INTEGER := 6;
	CONSTANT SERV_REQ       : INTEGER := 5;
	CONSTANT BROAD_COM      : INTEGER := 4;
	CONSTANT SUBSCR_BUSY    : INTEGER := 3;
	CONSTANT SUBSCR_ERR     : INTEGER := 2;
	CONSTANT BUS_CONTROL    : INTEGER := 1;
	CONSTANT TERMINAL_ERR   : INTEGER := 0;
	
	
	

	
	

END milstd_1553_pkg;
