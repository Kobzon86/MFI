LIBRARY IEEE;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.STD_LOGIC_1164.ALL;
USE work.i2c_heater_pkg.ALL;


PACKAGE lcd_heater_pkg IS
                                           -- PCIE_CoreCLK_OUT
	CONSTANT CLKIN_FREQ_HZ     : INTEGER := 625_000_000;             --62_500_000;
	CONSTANT I2C_CLK_FREQ_HZ   : INTEGER := 100_000;
	CONSTANT PWM_CLKIN_FREQ_HZ : INTEGER := 625_000;     --625_000;
	CONSTANT PWM_FREQ_HZ       : INTEGER := 200;
	CONSTANT PWM_MAX_VAL       : UNSIGNED( 15 DOWNTO 0 ) := x"1F40"; -- 8000 max pwm counter value

	CONSTANT AVM_ADDR_WIDTH    : INTEGER := 8; 
	CONSTANT AVM_DATA_WIDTH    : INTEGER := 32;
	CONSTANT AVCFG_ADDR_WIDTH  : INTEGER := 3;

	
	CONSTANT TERM1_I2C_ADDR    : STD_LOGIC_VECTOR( I2C_ADDR_WIDTH - 1 DOWNTO 0 ) := "1001000";  --DD1
	CONSTANT TERM2_I2C_ADDR    : STD_LOGIC_VECTOR( I2C_ADDR_WIDTH - 1 DOWNTO 0 ) := "1001001";  --DD2
	
	---------------- I2C TERMO SENSOR REGISTERS  ---------------------	
	CONSTANT I2CTERMO_TEMPER_ADDR   : STD_LOGIC_VECTOR( 7 DOWNTO 0 ) := x"00";	
	CONSTANT I2CTERMO_CFGREG_ADDR   : STD_LOGIC_VECTOR( 7 DOWNTO 0 ) := x"01";	
	CONSTANT I2CTERMO_HISTER_ADDR   : STD_LOGIC_VECTOR( 7 DOWNTO 0 ) := x"02";	
	CONSTANT I2CTERMO_OVTEMP_ADDR   : STD_LOGIC_VECTOR( 7 DOWNTO 0 ) := x"03";		
	
	
	----------------- Start timer interval ---------------------------
	CONSTANT TIMER_100MS        : STD_LOGIC_VECTOR( 19 DOWNTO 0 ) := STD_LOGIC_VECTOR( TO_UNSIGNED( 62500, 20 ) ); -- timer clock freq = 625000 Hz
	--CONSTANT TIMER_100MS        : STD_LOGIC_VECTOR( 19 DOWNTO 0 ) := STD_LOGIC_VECTOR( TO_UNSIGNED( 80000, 20 ) ); -- timer clock freq = 625000 Hz
	---------------- DEBUG ONLY ------------------------
	CONSTANT TIMER_1MS        : STD_LOGIC_VECTOR( 19 DOWNTO 0 ) := STD_LOGIC_VECTOR( TO_UNSIGNED( 625, 20 ) ); -- timer clock freq = 625000 Hz
	--CONSTANT TIMER_1MS        : STD_LOGIC_VECTOR( 19 DOWNTO 0 ) := STD_LOGIC_VECTOR( TO_UNSIGNED( 800, 20 ) ); -- timer clock freq = 625000 Hz
	
	------------------ LCD_Heater REGISTERS --------------------
	CONSTANT CONFIG_REG_ADDR    : INTEGER := 0;
	CONSTANT INTMASK_REG_ADDR   : INTEGER := 1;
	CONSTANT INTFLAG_REG_ADDR   : INTEGER := 2;
	
	------------------- CONFIG_REG BITS --------------
	CONSTANT TEMPER_H           : INTEGER := 8;
	CONSTANT TEMPER_L           : INTEGER := 1;
	CONSTANT HEATER_EN          : INTEGER := 0;
	
	------------------- INTFLAG_REG BITS -----------------
	CONSTANT SIGN_ERR_H         : INTEGER := 11;
	CONSTANT SIGN_ERR_L         : INTEGER := 10;
	CONSTANT TEMP_H             : INTEGER := 9;
	CONSTANT TEMP_L             : INTEGER := 3;
	CONSTANT TEMP2_ERR          : INTEGER := 2;
	CONSTANT TEMP1_ERR          : INTEGER := 1;
	CONSTANT PWM_ON             : INTEGER := 0;
	
	CONSTANT CLRBIT_H           : INTEGER := 2;
	CONSTANT CLRBIT_L           : INTEGER := 0;

	--CONSTANT SENSOR_ERROR_TEMPER : SIGNED( 6 DOWNTO 0 ) := TO_SIGNED( 10, 7 );  -- 10 degrees Celsius	
	
END lcd_heater_pkg;	
	
	
