LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;


PACKAGE i2c_swap_a429_pkg IS
	
		-------------- Avalon-MM width ----------------
	CONSTANT AVM_ADDR_WIDTH    : INTEGER := 20;
	CONSTANT AVM_DATA_WIDTH    : INTEGER := 32; 
	CONSTANT AVCFG_ADDR_WIDTH  : INTEGER := 4;
	
	CONSTANT FIFO_DATAWIDTH    : INTEGER := AVM_DATA_WIDTH;	
	CONSTANT FIFO_USEDWIDTH    : INTEGER := 10;
	CONSTANT FIFO_WORDNUM      : INTEGER := 1023;
	

	
	----------- A429RX Buffers Address Map ------------------------
	------------ A429 RxFIFO buffer address in file mode -------------
	CONSTANT A429RX_BUFF_ADDR    : UNSIGNED( AVM_ADDR_WIDTH - 1 DOWNTO 0 ) := resize( x"0000_0000"/4, AVM_ADDR_WIDTH );
	CONSTANT RXFIFO_OFFSET       : UNSIGNED( ( AVM_ADDR_WIDTH - 1 ) DOWNTO 0 ) := TO_UNSIGNED( 256, AVM_ADDR_WIDTH ); -- in ARINC429 Words  
	CONSTANT A429RX_FIFO_ADDR    : UNSIGNED( AVM_ADDR_WIDTH - 1 DOWNTO 0 ) := A429RX_BUFF_ADDR + RXFIFO_OFFSET;
	
	CONSTANT A429RX_CONFREG_ADDR : UNSIGNED( AVM_ADDR_WIDTH - 1 DOWNTO 0 ) := A429RX_BUFF_ADDR + resize( x"0000_4000"/4, AVM_ADDR_WIDTH );
	CONSTANT A429RX_INTREG_ADDR  : UNSIGNED( AVM_ADDR_WIDTH - 1 DOWNTO 0 ) := A429RX_CONFREG_ADDR + resize( x"0000_0008"/4, AVM_ADDR_WIDTH );  
	CONSTANT A429RX_BUFF_LEN     : UNSIGNED( AVM_ADDR_WIDTH - 1 DOWNTO 0 ) := TO_UNSIGNED( 768, AVM_ADDR_WIDTH );
	
-- 	CONSTANT A429RX_BUFF_ADDR_CHSTEP : UNSIGNED( AVM_ADDR_WIDTH - 1 DOWNTO 0 ) := resize( x"0001_0000"/4, AVM_ADDR_WIDTH );
	
	---------- A429RX0 CONFIG_REG Mapping -----------------
	CONSTANT CPU_BUFF_BUSY        : INTEGER := 26;
	CONSTANT ADDR_NROL            : INTEGER := 7;
	
	---------- A429RX0 INTFLAG_REG Mapping -----------------
	CONSTANT FPGA_BUFF_BUSY       : INTEGER := 26;
	CONSTANT RXWRD_AVAIL_H        : INTEGER := 25;
	CONSTANT RXWRD_AVAIL_L        : INTEGER := 16;
	CONSTANT RD_PTR_H             : INTEGER := 15;
	CONSTANT RD_PTR_L             : INTEGER := 6;
	
	
	
	------------ A429TX buffers Address Map ---------------------
	CONSTANT A429TX_BUFF_ADDR    : UNSIGNED( AVM_ADDR_WIDTH - 1 DOWNTO 0 ) := resize( x"0010_0000"/4, AVM_ADDR_WIDTH );
	CONSTANT A429TX_BUFF_LEN     : UNSIGNED( AVM_ADDR_WIDTH - 1 DOWNTO 0 ) := TO_UNSIGNED( 512, AVM_ADDR_WIDTH );
	CONSTANT A429TX_CONFREG_ADDR : UNSIGNED( AVM_ADDR_WIDTH - 1 DOWNTO 0 ) := A429TX_BUFF_ADDR + resize(x"0000_4000"/4, AVM_ADDR_WIDTH );
	CONSTANT A429TX_INTREG_ADDR  : UNSIGNED( AVM_ADDR_WIDTH - 1 DOWNTO 0 ) := A429TX_CONFREG_ADDR + resize( x"0000_0008"/4, AVM_ADDR_WIDTH );
 	
 		
	-------------- A429TX0 INTFLAG_REG Mapping ----------
	CONSTANT TX_FREESPACE_H    : INTEGER := 25;
	CONSTANT TX_FREESPACE_L    : INTEGER := 16;
	CONSTANT WR_PTR_H          : INTEGER := 15;
	CONSTANT WR_PTR_L          : INTEGER := 6;
	
	
	----------- I2C Buffers -----------------------------
	CONSTANT I2C_BUFF_ADDR     : UNSIGNED( AVM_ADDR_WIDTH - 1 DOWNTO 0 ) := resize( x"0020_0000"/4, AVM_ADDR_WIDTH );
--	CONSTANT I2C_TXBUFF_OFFSET : UNSIGNED( AVM_ADDR_WIDTH - 1 DOWNTO 0 ) := TO_UNSIGNED( 16, AVM_ADDR_WIDTH );
	CONSTANT I2C_TXBUFF_ADDR   : UNSIGNED( AVM_ADDR_WIDTH - 1 DOWNTO 0 ) := resize( x"0020_0040"/4, AVM_ADDR_WIDTH );  --I2C_BUFF_ADDR + I2C_TXBUFF_OFFSET;
	CONSTANT I2C_TXBUF_LEN     : UNSIGNED( AVM_ADDR_WIDTH - 1 DOWNTO 0 ) := TO_UNSIGNED( 16, AVM_ADDR_WIDTH );
	CONSTANT I2C_NIOS_BUFF_STARTADDR : UNSIGNED( AVM_ADDR_WIDTH - 1 DOWNTO 0 ) := resize( x"0021_0000"/4, AVM_ADDR_WIDTH );  --I2C_TXBUFF_ADDR + I2C_TXBUF_LEN;	
	--CONSTANT I2C_SWAP_DATA_LEN : UNSIGNED( ( RXWRD_AVAIL_H - RXWRD_AVAIL_L ) DOWNTO 0 ) := TO_UNSIGNED( 16, RXWRD_AVAIL_H - RXWRD_AVAIL_L + 1 );  
	CONSTANT I2C_SWAP_DATA_LEN : UNSIGNED( ( RXWRD_AVAIL_H - RXWRD_AVAIL_L ) DOWNTO 0 ) := TO_UNSIGNED( 16, RXWRD_AVAIL_H - RXWRD_AVAIL_L + 1 );  
	
	CONSTANT I2C_CONFREG_ADDR : UNSIGNED( AVM_ADDR_WIDTH - 1 DOWNTO 0 ) := I2C_BUFF_ADDR + resize(x"0000_4000"/4 ,AVM_ADDR_WIDTH );
	CONSTANT I2C_INTREG_ADDR  : UNSIGNED( AVM_ADDR_WIDTH - 1 DOWNTO 0 ) := I2C_CONFREG_ADDR + resize( x"0000_0008"/4, AVM_ADDR_WIDTH );
	
	
	
	---------- I2C INTFLAG_REG Mapping ----------------
	CONSTANT FPGA_RXBUFF_BUSY  : INTEGER := 26;
	CONSTANT FPGA_TXBUFF_BUSY  : INTEGER := 25;
	CONSTANT I2C_NEWDATA       : INTEGER := 0;
	
	------------ Internal Config Registers ----------------
	CONSTANT CONFIG_REG_ADDR     : INTEGER := 0;
	CONSTANT INTMASK_REG_ADDR    : INTEGER := 1;
	CONSTANT INTFLAG_REG_ADDR    : INTEGER := 2;


	
	--------------- CONFIG_REG BITS -------------------------------
	CONSTANT SWAP_EN             : INTEGER := 0;
	CONSTANT A429_CHAN_LB        : INTEGER := 1; -- select ARINC429 channel to swap data with I2C
	CONSTANT A429_CHAN_HB        : INTEGER := 5; -- select ARINC429 channel to swap data with I2C
	--CONSTANT I2C_FREQ_LB        : INTEGER := 1; -- 00 = 100 kHz, 01 = 50 kHz,
	--CONSTANT I2C_FREQ_HB        : INTEGER := 2; -- 10 = 25 kHz, 11 = 12.5 kHz
	--CONSTANT CPU_TXBUFF_BUSY    : INTEGER := 25;
	--CONSTANT CPU_RXBUFF_BUSY    : INTEGER := 26;
	
	
	
	
END i2c_swap_a429_pkg;	


	                     
	                     
	                     
